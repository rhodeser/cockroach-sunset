// n3_if_core.v - Digilent Nexys 3 board peripheral interface for ECE 544
//
// Copyright Copyright Roy Kravitz, Portland State University 2013, 2014, 2015
//
// Ported from the S3E Starter Board Interface by Roy Kravitz. Includes a simple 
// 8-bit interrupt controller for the PicoBlaze. The interrupt controller was derived
// from the simple interrupt controller from Opencores.org.  The two interrupt sources 
// are a 1ms clock tick used for debouncing the pushbuttons and switches and the rotary encoder event
// signal generated by the rotary_filter() module
//
// NOTES:
// ------
//	o	THIS INTERFACE REQUIRES THAT A DIGILENT PMODCLP (2 x 16 PARALLEL INTERFACE)
//		AND A PmodENC (ROTARY ENCODER WITH PUSHBUTTON AND SLIDE SWITCH) BE INSERTED
//		IN TWO OF THE PMOD EXPANSION CONNECTORS ON THE NEXYS 3.  THERE IS NO SIMPLE
//		WAY TO CHECK IF THE PERIPHERALS ARE INSERTED BO CAVEAT EMPTOR.
//
//	o	THIS VERSION OF THE INTERFACE CREATES AN 8-BIT INTERFACE TO THE PmodCLP. 
//		INITIALIZATION TIMING IS BASED ON A SAMSUNG KS0062U LCD CONTROLLER
//
//	o	THIS VERSION OF THE PROGRAM ONLY SUPPORTS THE LOW ORDER 4 SLIDE SWITCHES ON THE
//		NEXYS 3.  THIS IS DONE TO MAINTAIN BACKWARDS COMPATIBILITY WITH THE S3E STARTER
//		BOARD IMPLEMENTATION OF THE INTERFACE.  THE UPPER 4 SWITCHES AND TH SLIDE SWITCH
//		ON THE PmodENC CAN BE USED BY ADDING A GPIO PERIPHERAL TO YOUR XPS PROJECT	
//
// Created By:	Roy Kravitz
// Date:		13-March-2013
// Version:		1.0
//
// Description:
// ------------
// This module provides an interface to the Nexys 3 buttons, switches, and LEDs and to
// a PmodCLP and a PmodENC connected to 3 (PmodCLP uses two) Pmod expansion ports on
// the Nexys 3.  This design uses a Xilinx PicoBlaze to perform four distinct functions:
//	o 	pushbutton and switch debouncing -   The module debounces BTN_North, BTN_West and
// 		BTN_East and the rotary switch pushbuttons.  BTN_South is used as an FPGA reset signal
// 		in the Nexys 3 description file for the EDK so is not available for
// 		general use.   The module also debounces the lower 4 slide switches on the board.  
// 		Debounced buttons  and switches are:
//	 		db_btn_sw[7] - rotary_press (from the PmodENC)
//  		db_btn_sw[6] - btn_north (btnu in Nexys 3 documentation)
//  		db_btn_sw[5] - btn_east (btnl in Nexys 3 documentation)
//   		db_btn_sw[4] - btn_west (btnr in Nexys 3 documentation)
//			db_btn_sw[3] - slide switch 3
//			db_btn_sw[2] - slide switch 2 
//			db_btn_sw[1] - slide switch 1
//			db_btn_sw[0] - slide switch 0 (right most)
//
//	o	leds_out - The leds on the S3E board can be set by writing to the led_reg.
//
//	o	rotary encoder -  The rotary encoder delivers a 16-bit rotary_value[] register 
// 		that increments (decrements) every time the rotary encoder is moved to the
// 		right (left).  The rotary encoder is controlled by an 8-bit rotary_ctl[] input vector
//		with the following bits:
//			rotary_ctl[7]   = set the rotary_value to 0 when the signal is pulsed (0->1->0)
//			rotary_ctl[6]   = set the encoder increment value to rotary_ctl[3:0] when pulsed
//			rotary_ctl[5]   = reserved
//			rotary_ctl[4]   = set to limit the encoder values to >= 0  (no negative values)
//							  written when rotary_ctl[6] is pulsed.    
//			rotary_ctl[3:0] = increment/decrement interval for rotary_value[].  (default increment is 1)  
//
//			rotary_count_lo = least significant byte of rotary encoder count
//			rotary_count_hi = most significant byte of rotary encoder count
//			rotary_status   = returns the status of the rotary encoder control.  rotary_status[7] is a 'busy' flag
//							  which will be asserted high when the rotary encoder is busy.  rotary_status[6] is the
//							  'self test' flag.  It is asserted high while the s3 interface is doing its
//							  self test and deasserted when the self test is complete
//
//	o	lcd display - The LCD display on the PmodCLP is managed by the PicoBlaze software. An external
//		CPU (such as a microblaze or picoblaze) puts characters on the display and executes
//		display commands through three registers:
//			lcd_cmd - 	contains the LCD command.  when lcd_cmd[7] is toggled the cmd in lcd_cmd[4:0]
//						is translated and passed to the LCD display controller.
//			lcd_data -	contains the LCD data (character or display address)
//			lcd_status -returns the status of the LCD control.  At this point only
//						lcd_status[7] is used.  This bit is a 'busy' bit which will
//						be asserted high when the LCD display is busy.	
//	
// ***NOTE:  MODIFIED TO MAKE LCD_D AN OUTPUT - TAKES AWAY CAPABILITY OF READING *****
// ********  CHARACTER INFORMATION FROM THE LCD DISPLAY (NOT MUCH OF A LOSS)     *****
//////////////////////////////////////////////////////////////////////////////////////

module n3_if_core (
	// Nexys 3, PmodCLP and PmodENC interface
	// pushbuttons, switches and LEDs are on the Nexys 3.  Rotaty encoder and display
	// are provided with Digilent Pmods
	input				btn_west, btn_east,			// pushbutton inputs - left and right
	input				btn_north, rotary_press,	// pushbutton inputs - top and rotary_press
	input	[3:0]		sw,							// switch inputs
	input 				rotary_a, rotary_b, 		// rotary encoder inputs
	output	[7:0]		leds_out,					// led outputs
	
	// PmodCLP interface
	output				lcd_rs,						// LCD register select (1 = data)
						lcd_rw,						// LCD read/write (1 = read)
						lcd_e,						// LCD enable (1 = enable command)
	output	[7:0]		lcd_d,						// LCD data 
	
	// 1ms debounce clock - can be used w/ chipscope or for debug or for a timing signal
	output reg			db_clk,	
	
	// External CPU interface
	// Assumes that the inputs are instantiated as registers by the embedded CPU and 
	// are external to this module	
	
	// pushbuttons, switches and LEDs (Nexys 3)
	output	[7:0]		db_btn_sw,					// Debounced pushbuttons and switches
	input	[7:0]		leds_in,					// LED input values
	
	// rotary encoder (PmodENC)
	input	[7:0]		rotary_ctl,					// Rotary encoder control 
	output	[7:0]		rotary_count_lo,			// Rotary encoder count bits[7:0]
						rotary_count_hi,			// Rotary encoder count bits[15:8]
						rotary_status,				// Rotary encoder status
						
	// 16 x 2 LCD (PmodCLP)
	input	[7:0]		lcd_cmd,					// LCD command register
						lcd_data,					// LCD data register						
	output	[7:0]		lcd_status,					// LCD controller status		
	
	// System inputs
	input 				sysclk,            			// system clock
	input				sysreset					// system reset signal - asserted high to reset
);

	// I/O address ranges
	parameter  PBIF_START_ADDR = 8'd00,
	 	       PBIF_END_ADDR   = 8'd07,
	 	       PIC_START_ADDR  = 8'd08,
	 	       PIC_END_ADDR	   = 8'd15;


	
	//  declare internal variables
	
	// internal interface to/from the embedded Picoblaze in this s3e interface module
	wire	[7:0] 		port_id;
	wire   				write_strobe;
	wire   				read_strobe;
	wire	[7:0] 		out_port;
	wire	[7:0] 		in_port;
	wire	[9:0] 		address;
	wire	[17:0] 		instruction;
	wire				bram_enable;
	wire				rdl;
	wire				interrupt;
	wire				interrupt_ack;
	wire				kcpsm6_sleep;
	assign kcpsm6_sleep = 1'b0;
	
	wire				kcpsm6_reset; 
	assign kcpsm6_reset = rdl | sysreset;
	
	wire	[7:0]		btn_sw_in;					// buttons and switches input to picoblaze
	assign btn_sw_in = {rotary_press, btn_north, btn_east, btn_west, sw[3], sw[2], sw[1], sw[0]};
	
	wire				rotary_event;				// rotary encoder event - used as interrupt to picoblaze
	wire				rotary_left;				// rotary encoder direction - 1 says motion was to the left
	wire				db_rot_pbtn;				// debounced rotary pushbutton 
	assign db_rot_pbtn = db_btn_sw[7];				// This is bit 7 of the debounced button/switch register
	
	wire	[7:0]		lcd_ctl;					// LCD control signals driven by the picoblaze
	assign lcd_rs = lcd_ctl[2];
	assign lcd_rw = lcd_ctl[1];
	assign lcd_e = lcd_ctl[0];
	
	wire	[7:0]		lcd_dbus;					// LCD data bus driven by the picoblaze
	assign lcd_d = lcd_dbus;
	
	wire	[7:0]		rot_lcd_inputs;				// Rotary encoder and LCD inputs to picoblaze
	assign rot_lcd_inputs = {4'b0, 1'b0, db_rot_pbtn, rotary_event, rotary_left};
	
	// I/O interface enables
	wire				en_pic, en_pbif;			// enables for interrupt controller and PicoBlaze interface
	assign en_pic = (port_id >= PIC_START_ADDR) && (port_id <= PIC_END_ADDR);
	assign en_pbif = (port_id >= PBIF_START_ADDR) && (port_id <= PBIF_END_ADDR);
	
	// output buses from each of the I/O modules
	wire	[7:0]		pic_in_port, pbif_in_port;
	
	
	// instantiate the N3IF Ppcoblaze and its Program ROM
	kcpsm6 #(
		.interrupt_vector	(12'h3FF),
		.scratch_pad_memory_size(64),
		.hwbuild		(8'h00))
	N3IFCPU (
		.address 		(address),
		.instruction 	(instruction),
		.bram_enable 	(bram_enable),
		.port_id 		(port_id),
		.write_strobe 	(write_strobe),
		.k_write_strobe (),				// Constant Optimized writes are not used in this implementation
		.out_port 		(out_port),
		.read_strobe 	(read_strobe),
		.in_port 		(in_port),
		.interrupt 		(interrupt),
		.interrupt_ack 	(interrupt_ack),
		.reset 			(kcpsm6_reset),
		.sleep			(kcpsm6_sleep),
		.clk 			(sysclk)
); 

	// instantiate the firmware BRAM
	n3ifpgm #(
		.C_FAMILY		   ("S6"), 
		.C_RAM_SIZE_KWORDS	(1),
		.C_JTAG_LOADER_ENABLE	(1)) 
	N3IFPGM ( 
		.rdl 			(rdl),
		.enable 		(bram_enable),
		.address 		(address),
		.instruction 	(instruction),
		.clk 			(sysclk));
	
	// instantiate the interrupt controller
	pblaze_simple_pic 	PIC (
		.Wr_Strobe(write_strobe),
		.Rd_Strobe(read_strobe),
		.AddrIn(port_id),
		.DataIn(out_port),
		.DataOut(pic_in_port),
		.Int_in({6'b000000, rotary_event, db_clk}),
		.Int(interrupt),
		.Int_ack(interrupt_ack),	
		.enable(en_pic),
		.reset(sysreset),
		.clk(sysclk)
 	);
		
	// instantiate the rotary encoder filter
	// module is included in this file
	rotary_filter	RF (
		.rotary_a(rotary_a),
		.rotary_b(rotary_b),	
		.rotary_event(rotary_event),
		.rotary_left(rotary_left),				
		.clk(sysclk)
	);
	
	// instantiate the interface to the s3eif picoblaze
	pblaze_if  PBIF (
		// interface to/from the Picoblaze
		.Wr_Strobe(write_strobe),		// Write strobe - asserted to write I/O data
		.Rd_Strobe(read_strobe),		// Read strobe - asserted to read I/O data
		.AddrIn(port_id),				// I/O port address
		.DataIn(out_port),				// Data to be written to I/O register
		.DataOut(pbif_in_port),			// I/O register data to picoblaze
    	
    	
		// interface to the external CPU	
		.btn_sw_in(btn_sw_in),				// (I) buttons and switches from S3E board
		.leds_in(leds_in),					// (I) led contents to display
		.rotary_ctl(rotary_ctl),			// (I) rotary control register
		.rot_lcd_inputs(rot_lcd_inputs),	// (I) rotary encoder control and lcd data inputs
		.lcd_cmd(lcd_cmd),					// (I) LCD command register
		.lcd_data(lcd_data),				// (I) LCD data register
		
		.btn_sw_out(db_btn_sw),				// (O) debounced pushbuttons and switches
		.leds_out(leds_out),				// (O) led outputs
		.rotary_status(rotary_status),		// (O) rotary encoder status
		.rotary_count_lo(rotary_count_lo),	// (O) rotary count bits[7:0]
		.rotary_count_hi(rotary_count_hi),	// (O) rotary count bits[15:8]
		.lcd_status(lcd_status),			// (O) LCD status register
		.lcd_ctl(lcd_ctl),					// (O) LCD control signals
		.lcd_dbus(lcd_dbus),				// (O) LCD data bus

		.enable(en_pbif),		
   		.reset(sysreset),					// System reset
    	.clk(sysclk)						// 50Mhz clock signal
 	);
 
 	// Picoblaze input port data multiplexer
 	// defaults to Picoblaze interface except when PIC info is being written
	//assign in_port = en_pbif ? pbif_in_port : pic_in_port;
	assign in_port = en_pic ? pic_in_port : pbif_in_port;

 	// debounce clock - interrupt to s3 interface picoblaze
	parameter simulate = 0;
//	parameter simulate = 1;

    localparam debounce_cnt = simulate ? 21'd5          // debounce clock when simulating
                                       : 20'd0_100_000; // debounce count when running @ 100MHz on HW

	//internal registers	
	reg [19:0] db_count = 20'h00000;	//counter for debouncer
			
	always @(posedge sysclk)
	begin 
		if (db_count == debounce_cnt)begin
			db_clk <= 1;
			db_count <= 0;	//takes 1 mS to reach 100,000
		end
		else begin
			db_clk <= 0;
			db_count <= db_count + 1;
		end
	end	
	
		
endmodule
