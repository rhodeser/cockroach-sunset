//----------------------------------------------------------------------------
// user_logic.v - peripheral interface module for the Nexys 3 peripheral.
// the peripheral requires that a PmodCLP be connected to JA1 and JB1 and
// that a PmodENC be connected to the JC1 expansion connectors on the board
//----------------------------------------------------------------------------
//
// ***************************************************************************
// Copyright Roy Kravitz, Portland State University 2013, 2014, 2015
//
// Ported from the S3E Starter Board Interface by Roy Kravitz. Includes a simple 
// 8-bit interrupt controller for the PicoBlaze. The interrupt controller was derived
// from the simple interrupt controller from Opencores.org.  The two interrupt sources 
// are a 1ms clock tick used for debouncing the pushbuttons and switches and the rotary encoder event
// signal generated by the rotary_filter() module
//
// NOTES:
// ------
//	o	THIS INTERFACE REQUIRES THAT A DIGILENT PMODCLP (2 x 16 PARALLEL INTERFACE)
//		AND A PmodENC (ROTARY ENCODER WITH PUSHBUTTON AND SLIDE SWITCH) BE INSERTED
//		IN TWO OF THE PMOD EXPANSION CONNECTORS ON THE NEXYS 3.  THERE IS NO SIMPLE
//		WAY TO CHECK IF THE PERIPHERALS ARE INSERTED BO CAVEAT EMPTOR.
//
//	o	THIS VERSION OF THE INTERFACE CREATES AN 8-BIT INTERFACE TO THE PmodCLP. 
//		INITIALIZATION TIMING IS BASED ON A SAMSUNG KS0062U LCD CONTROLLER
//
//	o	THIS VERSION OF THE PROGRAM ONLY SUPPORTS THE LOW ORDER 4 SLIDE SWITCHES ON THE
//		NEXYS 3.  THIS IS DONE TO MAINTAIN BACKWARDS COMPATIBILITY WITH THE S3E STARTER
//		BOARD IMPLEMENTATION OF THE INTERFACE.  THE UPPER 4 SWITCHES AND TH SLIDE SWITCH
//		ON THE PmodENC CAN BE USED BY ADDING A GPIO PERIPHERAL TO YOUR XPS PROJECT	
//
// Created By:	Roy Kravitz
// Date:		13-March-2013
// Version:		1.0
//
// ***************************************************************************

// ***************************************************************************
// ** Copyright (c) 1995-2012 Xilinx, Inc.  All rights reserved.            **
// **                                                                       **
// ** Xilinx, Inc.                                                          **
// ** XILINX IS PROVIDING THIS DESIGN, CODE, OR INFORMATION "AS IS"         **
// ** AS A COURTESY TO YOU, SOLELY FOR USE IN DEVELOPING PROGRAMS AND       **
// ** SOLUTIONS FOR XILINX DEVICES.  BY PROVIDING THIS DESIGN, CODE,        **
// ** OR INFORMATION AS ONE POSSIBLE IMPLEMENTATION OF THIS FEATURE,        **
// ** APPLICATION OR STANDARD, XILINX IS MAKING NO REPRESENTATION           **
// ** THAT THIS IMPLEMENTATION IS FREE FROM ANY CLAIMS OF INFRINGEMENT,     **
// ** AND YOU ARE RESPONSIBLE FOR OBTAINING ANY RIGHTS YOU MAY REQUIRE      **
// ** FOR YOUR IMPLEMENTATION.  XILINX EXPRESSLY DISCLAIMS ANY              **
// ** WARRANTY WHATSOEVER WITH RESPECT TO THE ADEQUACY OF THE               **
// ** IMPLEMENTATION, INCLUDING BUT NOT LIMITED TO ANY WARRANTIES OR        **
// ** REPRESENTATIONS THAT THIS IMPLEMENTATION IS FREE FROM CLAIMS OF       **
// ** INFRINGEMENT, IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS       **
// ** FOR A PARTICULAR PURPOSE.                                             **
// **                                                                       **
// ***************************************************************************
//
//----------------------------------------------------------------------------
// Filename:          user_logic.v
// Version:           1.00.a
// Description:       User logic module.
// Date:              Thu Mar 14 06:09:39 2013 (by Create and Import Peripheral Wizard)
// Verilog Standard:  Verilog-2001
//----------------------------------------------------------------------------
// Naming Conventions:
//   active low signals:                    "*_n"
//   clock signals:                         "clk", "clk_div#", "clk_#x"
//   reset signals:                         "rst", "rst_n"
//   generics:                              "C_*"
//   user defined types:                    "*_TYPE"
//   state machine next state:              "*_ns"
//   state machine current state:           "*_cs"
//   combinatorial signals:                 "*_com"
//   pipelined or register delay signals:   "*_d#"
//   counter signals:                       "*cnt*"
//   clock enable signals:                  "*_ce"
//   internal version of output port:       "*_i"
//   device pins:                           "*_pin"
//   ports:                                 "- Names begin with Uppercase"
//   processes:                             "*_PROCESS"
//   component instantiations:              "<ENTITY_>I_<#|FUNC>"
//----------------------------------------------------------------------------

module user_logic
(
  // -- ADD USER PORTS BELOW THIS LINE ---------------
	btn_west,
	btn_east,
	btn_north,
	rotary_press,
	sw,
	rotary_a,
	rotary_b,
	leds_out,
	lcd_rs,
	lcd_rw,
	lcd_e,
	lcd_d,
	db_clk,	
  // -- ADD USER PORTS ABOVE THIS LINE ---------------

  // -- DO NOT EDIT BELOW THIS LINE ------------------
  // -- Bus protocol ports, do not add to or delete 
	Bus2IP_Clk,                     // Bus to IP clock
	Bus2IP_Reset,                   // Bus to IP reset
	Bus2IP_Data,                    // Bus to IP data bus
	Bus2IP_BE,                      // Bus to IP byte enables
	Bus2IP_RdCE,                    // Bus to IP read chip enable
	Bus2IP_WrCE,                    // Bus to IP write chip enable
	IP2Bus_Data,                    // IP to Bus data bus
	IP2Bus_RdAck,                   // IP to Bus read transfer acknowledgement
	IP2Bus_WrAck,                   // IP to Bus write transfer acknowledgement
	IP2Bus_Error                    // IP to Bus error response
  // -- DO NOT EDIT ABOVE THIS LINE ------------------
); // user_logic

// -- ADD USER PARAMETERS BELOW THIS LINE ------------
// ***** NO USER PARAMETERS *****
// -- ADD USER PARAMETERS ABOVE THIS LINE ------------

// -- DO NOT EDIT BELOW THIS LINE --------------------
// -- Bus protocol parameters, do not add to or delete
parameter C_SLV_DWIDTH                   = 32;
parameter C_NUM_REG                      = 10;
// -- DO NOT EDIT ABOVE THIS LINE --------------------

// -- ADD USER PORTS BELOW THIS LINE -----------------
input									btn_west;		// Nexys 3 pushbutton inputs - left, right, and up
input									btn_east;
input									btn_north;
input									rotary_press;	// PmodENC rotary encoder pushbutton
input	[3:0]							sw;				// Nexys 3 switch inputs
input 									rotary_a;		// PmodENC rotary encoder inputs
input									rotary_b;
output	[7:0]							leds_out;		// Nexys 3 LED outputs

output									lcd_rs;			// PmodCLP LCD register select (1 = data)
output									lcd_rw;			// PmosCLP LCD read/write (1 = read)
output									lcd_e;			// PmodCLP LCD enable (1 = enable command)
output	[7:0]							lcd_d;			// PmodCLP LCD data 
output									db_clk;			//1ms debounce clock - can be used for debug or slow clock
// -- ADD USER PORTS ABOVE THIS LINE -----------------

// -- DO NOT EDIT BELOW THIS LINE --------------------
// -- Bus protocol ports, do not add to or delete
input                                     Bus2IP_Clk;
input                                     Bus2IP_Reset;
input      [0 : C_SLV_DWIDTH-1]           Bus2IP_Data;
input      [0 : C_SLV_DWIDTH/8-1]         Bus2IP_BE;
input      [0 : C_NUM_REG-1]              Bus2IP_RdCE;
input      [0 : C_NUM_REG-1]              Bus2IP_WrCE;
output     [0 : C_SLV_DWIDTH-1]           IP2Bus_Data;
output                                    IP2Bus_RdAck;
output                                    IP2Bus_WrAck;
output                                    IP2Bus_Error;
// -- DO NOT EDIT ABOVE THIS LINE --------------------

//----------------------------------------------------------------------------
// Implementation
//----------------------------------------------------------------------------

  // --USER nets declarations added here, as needed for user logic
  wire		[7:0]							db_btn_sw;					// Debounced pushbuttons and switches
  wire		[7:0]							leds_in;					// LED input values
  wire		[7:0]							rotary_ctl;					// Rotary encoder control 
  wire		[7:0]							rotary_count_lo;			// Rotary encoder count bits[7:0]
  wire		[7:0]							rotary_count_hi;			// Rotary encoder count bits[15:8]
  wire		[7:0]							rotary_status;				// Rotary encoder status
  wire		[7:0]							lcd_cmd;					// LCD command register
  wire		[7:0]							lcd_data;					// LCD data register						
  wire		[7:0]							lcd_status;					// LCD controller status
  
  // Nets for user logic slave model s/w accessible register example
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg0;
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg1;
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg2;
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg3;
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg4;
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg5;
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg6;
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg7;
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg8;
  reg        [0 : C_SLV_DWIDTH-1]           slv_reg9;
  wire       [0 : 9]                        slv_reg_write_sel;
  wire       [0 : 9]                        slv_reg_read_sel;
  reg        [0 : C_SLV_DWIDTH-1]           slv_ip2bus_data;
  wire                                      slv_read_ack;
  wire                                      slv_write_ack;
  integer                                   byte_index, bit_index;

  // --USER logic implementation added here
  
  // instantiate the core peripheral
  n3_if_core N3IF (
	.btn_west(btn_west),
	.btn_east(btn_east),
	.btn_north(btn_north),
	.rotary_press(rotary_press),
	.sw(sw),
	.rotary_a(rotary_a),
	.rotary_b(rotary_b),
	.leds_out(leds_out),
	.lcd_rs(lcd_rs),
	.lcd_rw(lcd_rw),
	.lcd_e(lcd_e),
	.lcd_d(lcd_d),
	.db_clk(db_clk),	
	.db_btn_sw(db_btn_sw),
	.leds_in(leds_in),
	.rotary_ctl(rotary_ctl),
	.rotary_count_lo(rotary_count_lo),
	.rotary_count_hi(rotary_count_hi),
	.rotary_status(rotary_status),
	.lcd_cmd(lcd_cmd),
	.lcd_data(lcd_data),			
	.lcd_status(lcd_status),
	.sysclk(Bus2IP_Clk),
	.sysreset(Bus2IP_Reset)	
);

// Assign the slave registers based on their memory mapped address

// microblaze input registers (from periperal to microblaze)
always @* begin
	slv_reg0 = {24'h000000, db_btn_sw};
	slv_reg1 = {24'h000000, rotary_status};
	slv_reg2 = {24'h000000, rotary_count_lo}; 
	slv_reg3 = {24'h000000, rotary_count_hi};
	slv_reg4 = {24'h000000, lcd_status};
end // assign microblaze input registers

// microblaze output registers (from microblaze to peripheral)
assign leds_in = slv_reg5[24:31];
assign rotary_ctl = slv_reg6[24:31];
assign lcd_cmd = slv_reg7[24:31];
assign lcd_data = slv_reg8[24:31];

  // ------------------------------------------------------
  // Example code to read/write user logic slave model s/w accessible registers
  // 
  // Note:
  // The example code presented here is to show you one way of reading/writing
  // software accessible registers implemented in the user logic slave model.
  // Each bit of the Bus2IP_WrCE/Bus2IP_RdCE signals is configured to correspond
  // to one software accessible register by the top level template. For example,
  // if you have four 32 bit software accessible registers in the user logic,
  // you are basically operating on the following memory mapped registers:
  // 
  //    Bus2IP_WrCE/Bus2IP_RdCE   Memory Mapped Register
  //                     "1000"   C_BASEADDR + 0x0
  //                     "0100"   C_BASEADDR + 0x4
  //                     "0010"   C_BASEADDR + 0x8
  //                     "0001"   C_BASEADDR + 0xC
  // 
  // ------------------------------------------------------

  assign
    slv_reg_write_sel = Bus2IP_WrCE[0:9],
    slv_reg_read_sel  = Bus2IP_RdCE[0:9],
    slv_write_ack     = Bus2IP_WrCE[0] || Bus2IP_WrCE[1] || Bus2IP_WrCE[2] || Bus2IP_WrCE[3] || Bus2IP_WrCE[4] || Bus2IP_WrCE[5] || Bus2IP_WrCE[6] || Bus2IP_WrCE[7] || Bus2IP_WrCE[8] || Bus2IP_WrCE[9],
    slv_read_ack      = Bus2IP_RdCE[0] || Bus2IP_RdCE[1] || Bus2IP_RdCE[2] || Bus2IP_RdCE[3] || Bus2IP_RdCE[4] || Bus2IP_RdCE[5] || Bus2IP_RdCE[6] || Bus2IP_RdCE[7] || Bus2IP_RdCE[8] || Bus2IP_RdCE[9];

  // implement slave model register(s)
  always @( posedge Bus2IP_Clk )
    begin: SLAVE_REG_WRITE_PROC

      if ( Bus2IP_Reset == 1 )
        begin
		/* These registers are read-only and assigned by the n3_if_core
			slv_reg0 <= 0;
			slv_reg1 <= 0;
			slv_reg2 <= 0;
			slv_reg3 <= 0;
			slv_reg4 <= 0;
		*/
		
          slv_reg5 <= 0;
          slv_reg6 <= 0;
          slv_reg7 <= 0;
          slv_reg8 <= 0;
          slv_reg9 <= 0;
        end
      else
        case ( slv_reg_write_sel )
		/* These registers are read-only and assigned by the n3_if_core
          10'b1000000000 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg0[bit_index] <= Bus2IP_Data[bit_index];
          10'b0100000000 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg1[bit_index] <= Bus2IP_Data[bit_index];
          10'b0010000000 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg2[bit_index] <= Bus2IP_Data[bit_index];
          10'b0001000000 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg3[bit_index] <= Bus2IP_Data[bit_index];
          10'b0000100000 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg4[bit_index] <= Bus2IP_Data[bit_index];
		*/
		
          10'b0000010000 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg5[bit_index] <= Bus2IP_Data[bit_index];
          10'b0000001000 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg6[bit_index] <= Bus2IP_Data[bit_index];
          10'b0000000100 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg7[bit_index] <= Bus2IP_Data[bit_index];
          10'b0000000010 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg8[bit_index] <= Bus2IP_Data[bit_index];
						
          10'b0000000001 :
            for ( byte_index = 0; byte_index <= (C_SLV_DWIDTH/8)-1; byte_index = byte_index+1 )
              if ( Bus2IP_BE[byte_index] == 1 )
                for ( bit_index = byte_index*8; bit_index <= byte_index*8+7; bit_index = bit_index+1 )
                  slv_reg9[bit_index] <= Bus2IP_Data[bit_index];
			
          default : ;
        endcase

    end // SLAVE_REG_WRITE_PROC

  // implement slave model register read mux
  always @( slv_reg_read_sel or slv_reg0 or slv_reg1 or slv_reg2 or slv_reg3 or slv_reg4 or slv_reg5 or slv_reg6 or slv_reg7 or slv_reg8 or slv_reg9 )
    begin: SLAVE_REG_READ_PROC

      case ( slv_reg_read_sel )
        10'b1000000000 : slv_ip2bus_data <= slv_reg0;
        10'b0100000000 : slv_ip2bus_data <= slv_reg1;
        10'b0010000000 : slv_ip2bus_data <= slv_reg2;
        10'b0001000000 : slv_ip2bus_data <= slv_reg3;
        10'b0000100000 : slv_ip2bus_data <= slv_reg4;
        10'b0000010000 : slv_ip2bus_data <= slv_reg5;
        10'b0000001000 : slv_ip2bus_data <= slv_reg6;
        10'b0000000100 : slv_ip2bus_data <= slv_reg7;
        10'b0000000010 : slv_ip2bus_data <= slv_reg8;
        10'b0000000001 : slv_ip2bus_data <= slv_reg9;
        default : slv_ip2bus_data <= 0;
      endcase

    end // SLAVE_REG_READ_PROC

  // ------------------------------------------------------------
  // Example code to drive IP to Bus signals
  // ------------------------------------------------------------

  assign IP2Bus_Data    = slv_ip2bus_data;
  assign IP2Bus_WrAck   = slv_write_ack;
  assign IP2Bus_RdAck   = slv_read_ack;
  assign IP2Bus_Error   = 0;

endmodule
